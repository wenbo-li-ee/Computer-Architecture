VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_2rw_64x128_64
   CLASS BLOCK ;
   SIZE 535.54 BY 425.38 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.72 0.0 105.1 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.84 0.0 111.22 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.28 0.0 116.66 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.08 0.0 123.46 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  128.52 0.0 128.9 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.96 0.0 134.34 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.08 0.0 140.46 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  145.52 0.0 145.9 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  152.32 0.0 152.7 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 0.0 158.14 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 0.0 163.58 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.32 0.0 169.7 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  175.44 0.0 175.82 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.88 0.0 181.26 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 0.0 186.7 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  199.24 0.0 199.62 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.68 0.0 205.06 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 0.0 210.5 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.68 0.0 222.06 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 0.0 228.18 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.92 0.0 234.3 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  239.36 0.0 239.74 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.8 0.0 245.18 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  251.6 0.0 251.98 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 0.0 257.42 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 0.0 269.66 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 0.0 274.42 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 0.0 281.22 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 0.0 286.66 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  291.72 0.0 292.1 1.06 ;
      END
   END din0[32]
   PIN din0[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 0.0 298.22 1.06 ;
      END
   END din0[33]
   PIN din0[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  303.28 0.0 303.66 1.06 ;
      END
   END din0[34]
   PIN din0[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 0.0 310.46 1.06 ;
      END
   END din0[35]
   PIN din0[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  315.52 0.0 315.9 1.06 ;
      END
   END din0[36]
   PIN din0[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  320.96 0.0 321.34 1.06 ;
      END
   END din0[37]
   PIN din0[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  327.76 0.0 328.14 1.06 ;
      END
   END din0[38]
   PIN din0[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  333.2 0.0 333.58 1.06 ;
      END
   END din0[39]
   PIN din0[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  338.64 0.0 339.02 1.06 ;
      END
   END din0[40]
   PIN din0[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.08 0.0 344.46 1.06 ;
      END
   END din0[41]
   PIN din0[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  350.2 0.0 350.58 1.06 ;
      END
   END din0[42]
   PIN din0[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  355.64 0.0 356.02 1.06 ;
      END
   END din0[43]
   PIN din0[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  362.44 0.0 362.82 1.06 ;
      END
   END din0[44]
   PIN din0[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  367.88 0.0 368.26 1.06 ;
      END
   END din0[45]
   PIN din0[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  373.32 0.0 373.7 1.06 ;
      END
   END din0[46]
   PIN din0[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 0.0 379.82 1.06 ;
      END
   END din0[47]
   PIN din0[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  384.88 0.0 385.26 1.06 ;
      END
   END din0[48]
   PIN din0[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  391.68 0.0 392.06 1.06 ;
      END
   END din0[49]
   PIN din0[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  397.12 0.0 397.5 1.06 ;
      END
   END din0[50]
   PIN din0[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  402.56 0.0 402.94 1.06 ;
      END
   END din0[51]
   PIN din0[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  409.36 0.0 409.74 1.06 ;
      END
   END din0[52]
   PIN din0[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  414.8 0.0 415.18 1.06 ;
      END
   END din0[53]
   PIN din0[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  420.24 0.0 420.62 1.06 ;
      END
   END din0[54]
   PIN din0[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  426.36 0.0 426.74 1.06 ;
      END
   END din0[55]
   PIN din0[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  431.8 0.0 432.18 1.06 ;
      END
   END din0[56]
   PIN din0[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  438.6 0.0 438.98 1.06 ;
      END
   END din0[57]
   PIN din0[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  444.04 0.0 444.42 1.06 ;
      END
   END din0[58]
   PIN din0[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  449.48 0.0 449.86 1.06 ;
      END
   END din0[59]
   PIN din0[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  454.92 0.0 455.3 1.06 ;
      END
   END din0[60]
   PIN din0[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  461.04 0.0 461.42 1.06 ;
      END
   END din0[61]
   PIN din0[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  467.16 0.0 467.54 1.06 ;
      END
   END din0[62]
   PIN din0[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  473.28 0.0 473.66 1.06 ;
      END
   END din0[63]
   PIN din1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  51.68 424.32 52.06 425.38 ;
      END
   END din1[0]
   PIN din1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  58.48 424.32 58.86 425.38 ;
      END
   END din1[1]
   PIN din1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  64.6 424.32 64.98 425.38 ;
      END
   END din1[2]
   PIN din1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  70.04 424.32 70.42 425.38 ;
      END
   END din1[3]
   PIN din1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  75.48 424.32 75.86 425.38 ;
      END
   END din1[4]
   PIN din1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.92 424.32 81.3 425.38 ;
      END
   END din1[5]
   PIN din1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.72 424.32 88.1 425.38 ;
      END
   END din1[6]
   PIN din1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.16 424.32 93.54 425.38 ;
      END
   END din1[7]
   PIN din1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.6 424.32 98.98 425.38 ;
      END
   END din1[8]
   PIN din1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  105.4 424.32 105.78 425.38 ;
      END
   END din1[9]
   PIN din1[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.84 424.32 111.22 425.38 ;
      END
   END din1[10]
   PIN din1[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.96 424.32 117.34 425.38 ;
      END
   END din1[11]
   PIN din1[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  122.4 424.32 122.78 425.38 ;
      END
   END din1[12]
   PIN din1[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.84 424.32 128.22 425.38 ;
      END
   END din1[13]
   PIN din1[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.96 424.32 134.34 425.38 ;
      END
   END din1[14]
   PIN din1[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.08 424.32 140.46 425.38 ;
      END
   END din1[15]
   PIN din1[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  146.2 424.32 146.58 425.38 ;
      END
   END din1[16]
   PIN din1[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  151.64 424.32 152.02 425.38 ;
      END
   END din1[17]
   PIN din1[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.08 424.32 157.46 425.38 ;
      END
   END din1[18]
   PIN din1[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 424.32 163.58 425.38 ;
      END
   END din1[19]
   PIN din1[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.32 424.32 169.7 425.38 ;
      END
   END din1[20]
   PIN din1[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.76 424.32 175.14 425.38 ;
      END
   END din1[21]
   PIN din1[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 424.32 180.58 425.38 ;
      END
   END din1[22]
   PIN din1[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  187.0 424.32 187.38 425.38 ;
      END
   END din1[23]
   PIN din1[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 424.32 192.82 425.38 ;
      END
   END din1[24]
   PIN din1[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  198.56 424.32 198.94 425.38 ;
      END
   END din1[25]
   PIN din1[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 424.32 204.38 425.38 ;
      END
   END din1[26]
   PIN din1[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  209.44 424.32 209.82 425.38 ;
      END
   END din1[27]
   PIN din1[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 424.32 216.62 425.38 ;
      END
   END din1[28]
   PIN din1[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.68 424.32 222.06 425.38 ;
      END
   END din1[29]
   PIN din1[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 424.32 228.18 425.38 ;
      END
   END din1[30]
   PIN din1[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 424.32 232.94 425.38 ;
      END
   END din1[31]
   PIN din1[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 424.32 239.06 425.38 ;
      END
   END din1[32]
   PIN din1[33]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  245.48 424.32 245.86 425.38 ;
      END
   END din1[33]
   PIN din1[34]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 424.32 251.3 425.38 ;
      END
   END din1[34]
   PIN din1[35]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  256.36 424.32 256.74 425.38 ;
      END
   END din1[35]
   PIN din1[36]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.8 424.32 262.18 425.38 ;
      END
   END din1[36]
   PIN din1[37]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  268.6 424.32 268.98 425.38 ;
      END
   END din1[37]
   PIN din1[38]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.72 424.32 275.1 425.38 ;
      END
   END din1[38]
   PIN din1[39]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  280.16 424.32 280.54 425.38 ;
      END
   END din1[39]
   PIN din1[40]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  285.6 424.32 285.98 425.38 ;
      END
   END din1[40]
   PIN din1[41]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 424.32 291.42 425.38 ;
      END
   END din1[41]
   PIN din1[42]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 424.32 298.22 425.38 ;
      END
   END din1[42]
   PIN din1[43]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  303.96 424.32 304.34 425.38 ;
      END
   END din1[43]
   PIN din1[44]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 424.32 309.78 425.38 ;
      END
   END din1[44]
   PIN din1[45]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  314.84 424.32 315.22 425.38 ;
      END
   END din1[45]
   PIN din1[46]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  320.28 424.32 320.66 425.38 ;
      END
   END din1[46]
   PIN din1[47]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  327.08 424.32 327.46 425.38 ;
      END
   END din1[47]
   PIN din1[48]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  332.52 424.32 332.9 425.38 ;
      END
   END din1[48]
   PIN din1[49]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  337.96 424.32 338.34 425.38 ;
      END
   END din1[49]
   PIN din1[50]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  344.76 424.32 345.14 425.38 ;
      END
   END din1[50]
   PIN din1[51]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  350.2 424.32 350.58 425.38 ;
      END
   END din1[51]
   PIN din1[52]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  356.32 424.32 356.7 425.38 ;
      END
   END din1[52]
   PIN din1[53]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  361.08 424.32 361.46 425.38 ;
      END
   END din1[53]
   PIN din1[54]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  367.2 424.32 367.58 425.38 ;
      END
   END din1[54]
   PIN din1[55]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  374.0 424.32 374.38 425.38 ;
      END
   END din1[55]
   PIN din1[56]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  379.44 424.32 379.82 425.38 ;
      END
   END din1[56]
   PIN din1[57]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  385.56 424.32 385.94 425.38 ;
      END
   END din1[57]
   PIN din1[58]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  391.0 424.32 391.38 425.38 ;
      END
   END din1[58]
   PIN din1[59]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  396.44 424.32 396.82 425.38 ;
      END
   END din1[59]
   PIN din1[60]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  402.56 424.32 402.94 425.38 ;
      END
   END din1[60]
   PIN din1[61]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  408.68 424.32 409.06 425.38 ;
      END
   END din1[61]
   PIN din1[62]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  414.12 424.32 414.5 425.38 ;
      END
   END din1[62]
   PIN din1[63]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  419.56 424.32 419.94 425.38 ;
      END
   END din1[63]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 121.72 1.06 122.1 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 131.24 1.06 131.62 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 137.36 1.06 137.74 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 143.48 1.06 143.86 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 150.28 1.06 150.66 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 158.44 1.06 158.82 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.88 1.06 164.26 ;
      END
   END addr0[6]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  437.92 0.0 438.3 1.06 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  444.72 0.0 445.1 1.06 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  439.28 0.0 439.66 1.06 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  439.96 0.0 440.34 1.06 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  440.64 0.0 441.02 1.06 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  442.0 0.0 442.38 1.06 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  441.32 0.0 441.7 1.06 ;
      END
   END addr1[6]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 21.08 1.06 21.46 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  534.48 391.0 535.54 391.38 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 30.6 1.06 30.98 ;
      END
   END web0
   PIN web1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  534.48 382.84 535.54 383.22 ;
      END
   END web1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  30.6 0.0 30.98 1.06 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  534.48 389.64 535.54 390.02 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.28 0.0 167.66 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 0.0 173.1 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.4 0.0 173.78 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 0.0 179.22 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 0.0 182.62 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.96 0.0 185.34 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.0 0.0 187.38 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 0.0 193.5 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.8 0.0 194.18 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.56 0.0 198.94 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  199.92 0.0 200.3 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 0.0 204.38 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 0.0 205.74 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.8 0.0 211.18 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 0.0 211.86 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 0.0 217.3 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 0.0 217.98 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 0.0 223.42 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 0.0 224.78 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 0.0 230.22 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 0.0 230.9 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.28 0.0 235.66 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  236.64 0.0 237.02 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 0.0 241.78 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.76 0.0 243.14 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 0.0 248.58 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 0.0 249.26 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  254.32 0.0 254.7 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.0 0.0 255.38 1.06 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  260.44 0.0 260.82 1.06 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.84 0.0 264.22 1.06 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.56 0.0 266.94 1.06 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  268.6 0.0 268.98 1.06 ;
      END
   END dout0[32]
   PIN dout0[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.68 0.0 273.06 1.06 ;
      END
   END dout0[33]
   PIN dout0[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  274.72 0.0 275.1 1.06 ;
      END
   END dout0[34]
   PIN dout0[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 0.0 278.5 1.06 ;
      END
   END dout0[35]
   PIN dout0[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.16 0.0 280.54 1.06 ;
      END
   END dout0[36]
   PIN dout0[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.24 0.0 284.62 1.06 ;
      END
   END dout0[37]
   PIN dout0[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.96 0.0 287.34 1.06 ;
      END
   END dout0[38]
   PIN dout0[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  292.4 0.0 292.78 1.06 ;
      END
   END dout0[39]
   PIN dout0[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  293.08 0.0 293.46 1.06 ;
      END
   END dout0[40]
   PIN dout0[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  298.52 0.0 298.9 1.06 ;
      END
   END dout0[41]
   PIN dout0[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  299.2 0.0 299.58 1.06 ;
      END
   END dout0[42]
   PIN dout0[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 0.0 305.02 1.06 ;
      END
   END dout0[43]
   PIN dout0[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  305.32 0.0 305.7 1.06 ;
      END
   END dout0[44]
   PIN dout0[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.76 0.0 311.14 1.06 ;
      END
   END dout0[45]
   PIN dout0[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  311.44 0.0 311.82 1.06 ;
      END
   END dout0[46]
   PIN dout0[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.88 0.0 317.26 1.06 ;
      END
   END dout0[47]
   PIN dout0[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 0.0 317.94 1.06 ;
      END
   END dout0[48]
   PIN dout0[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.0 0.0 323.38 1.06 ;
      END
   END dout0[49]
   PIN dout0[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.68 0.0 324.06 1.06 ;
      END
   END dout0[50]
   PIN dout0[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.12 0.0 329.5 1.06 ;
      END
   END dout0[51]
   PIN dout0[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 0.0 330.86 1.06 ;
      END
   END dout0[52]
   PIN dout0[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.24 0.0 335.62 1.06 ;
      END
   END dout0[53]
   PIN dout0[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  336.6 0.0 336.98 1.06 ;
      END
   END dout0[54]
   PIN dout0[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 0.0 341.74 1.06 ;
      END
   END dout0[55]
   PIN dout0[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.72 0.0 343.1 1.06 ;
      END
   END dout0[56]
   PIN dout0[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.16 0.0 348.54 1.06 ;
      END
   END dout0[57]
   PIN dout0[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.88 0.0 351.26 1.06 ;
      END
   END dout0[58]
   PIN dout0[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  353.6 0.0 353.98 1.06 ;
      END
   END dout0[59]
   PIN dout0[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  354.28 0.0 354.66 1.06 ;
      END
   END dout0[60]
   PIN dout0[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  359.72 0.0 360.1 1.06 ;
      END
   END dout0[61]
   PIN dout0[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  361.76 0.0 362.14 1.06 ;
      END
   END dout0[62]
   PIN dout0[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  368.56 0.0 368.94 1.06 ;
      END
   END dout0[63]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.6 424.32 166.98 425.38 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.72 424.32 173.1 425.38 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 424.32 176.5 425.38 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.84 424.32 179.22 425.38 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 424.32 182.62 425.38 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 424.32 186.7 425.38 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.68 424.32 188.06 425.38 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.12 424.32 193.5 425.38 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.8 424.32 194.18 425.38 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.88 424.32 198.26 425.38 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  199.24 424.32 199.62 425.38 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  204.68 424.32 205.06 425.38 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.36 424.32 205.74 425.38 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 424.32 210.5 425.38 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.48 424.32 211.86 425.38 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.92 424.32 217.3 425.38 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.6 424.32 217.98 425.38 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  223.04 424.32 223.42 425.38 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 424.32 224.78 425.38 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  229.84 424.32 230.22 425.38 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 424.32 230.9 425.38 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.28 424.32 235.66 425.38 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  236.64 424.32 237.02 425.38 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  241.4 424.32 241.78 425.38 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  242.76 424.32 243.14 425.38 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 424.32 248.58 425.38 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.88 424.32 249.26 425.38 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  254.32 424.32 254.7 425.38 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 424.32 257.42 425.38 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  260.44 424.32 260.82 425.38 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.84 424.32 264.22 425.38 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  267.92 424.32 268.3 425.38 ;
      END
   END dout1[31]
   PIN dout1[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.96 424.32 270.34 425.38 ;
      END
   END dout1[32]
   PIN dout1[33]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 424.32 274.42 425.38 ;
      END
   END dout1[33]
   PIN dout1[34]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 424.32 276.46 425.38 ;
      END
   END dout1[34]
   PIN dout1[35]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.12 424.32 278.5 425.38 ;
      END
   END dout1[35]
   PIN dout1[36]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.84 424.32 281.22 425.38 ;
      END
   END dout1[36]
   PIN dout1[37]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 424.32 286.66 425.38 ;
      END
   END dout1[37]
   PIN dout1[38]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.96 424.32 287.34 425.38 ;
      END
   END dout1[38]
   PIN dout1[39]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  291.72 424.32 292.1 425.38 ;
      END
   END dout1[39]
   PIN dout1[40]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  293.08 424.32 293.46 425.38 ;
      END
   END dout1[40]
   PIN dout1[41]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  298.52 424.32 298.9 425.38 ;
      END
   END dout1[41]
   PIN dout1[42]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  299.2 424.32 299.58 425.38 ;
      END
   END dout1[42]
   PIN dout1[43]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 424.32 305.02 425.38 ;
      END
   END dout1[43]
   PIN dout1[44]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  305.32 424.32 305.7 425.38 ;
      END
   END dout1[44]
   PIN dout1[45]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  310.08 424.32 310.46 425.38 ;
      END
   END dout1[45]
   PIN dout1[46]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  311.44 424.32 311.82 425.38 ;
      END
   END dout1[46]
   PIN dout1[47]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.88 424.32 317.26 425.38 ;
      END
   END dout1[47]
   PIN dout1[48]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  317.56 424.32 317.94 425.38 ;
      END
   END dout1[48]
   PIN dout1[49]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.0 424.32 323.38 425.38 ;
      END
   END dout1[49]
   PIN dout1[50]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  323.68 424.32 324.06 425.38 ;
      END
   END dout1[50]
   PIN dout1[51]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  329.12 424.32 329.5 425.38 ;
      END
   END dout1[51]
   PIN dout1[52]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  330.48 424.32 330.86 425.38 ;
      END
   END dout1[52]
   PIN dout1[53]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.24 424.32 335.62 425.38 ;
      END
   END dout1[53]
   PIN dout1[54]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.92 424.32 336.3 425.38 ;
      END
   END dout1[54]
   PIN dout1[55]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  341.36 424.32 341.74 425.38 ;
      END
   END dout1[55]
   PIN dout1[56]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  342.04 424.32 342.42 425.38 ;
      END
   END dout1[56]
   PIN dout1[57]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  348.16 424.32 348.54 425.38 ;
      END
   END dout1[57]
   PIN dout1[58]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  350.88 424.32 351.26 425.38 ;
      END
   END dout1[58]
   PIN dout1[59]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  353.6 424.32 353.98 425.38 ;
      END
   END dout1[59]
   PIN dout1[60]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  357.0 424.32 357.38 425.38 ;
      END
   END dout1[60]
   PIN dout1[61]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  359.72 424.32 360.1 425.38 ;
      END
   END dout1[61]
   PIN dout1[62]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  361.76 424.32 362.14 425.38 ;
      END
   END dout1[62]
   PIN dout1[63]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  367.88 424.32 368.26 425.38 ;
      END
   END dout1[63]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  4.76 4.76 530.78 6.5 ;
         LAYER met4 ;
         RECT  4.76 4.76 6.5 420.62 ;
         LAYER met3 ;
         RECT  4.76 418.88 530.78 420.62 ;
         LAYER met4 ;
         RECT  529.04 4.76 530.78 420.62 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  532.44 1.36 534.18 424.02 ;
         LAYER met3 ;
         RECT  1.36 422.28 534.18 424.02 ;
         LAYER met4 ;
         RECT  1.36 1.36 3.1 424.02 ;
         LAYER met3 ;
         RECT  1.36 1.36 534.18 3.1 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 534.92 424.76 ;
   LAYER  met2 ;
      RECT  0.62 0.62 534.92 424.76 ;
   LAYER  met3 ;
      RECT  1.66 121.12 534.92 122.7 ;
      RECT  0.62 122.7 1.66 130.64 ;
      RECT  0.62 132.22 1.66 136.76 ;
      RECT  0.62 138.34 1.66 142.88 ;
      RECT  0.62 144.46 1.66 149.68 ;
      RECT  0.62 151.26 1.66 157.84 ;
      RECT  0.62 159.42 1.66 163.28 ;
      RECT  1.66 122.7 533.88 390.4 ;
      RECT  1.66 390.4 533.88 391.98 ;
      RECT  0.62 22.06 1.66 30.0 ;
      RECT  0.62 31.58 1.66 121.12 ;
      RECT  533.88 122.7 534.92 382.24 ;
      RECT  533.88 383.82 534.92 389.04 ;
      RECT  1.66 4.16 4.16 7.1 ;
      RECT  1.66 7.1 4.16 121.12 ;
      RECT  4.16 7.1 531.38 121.12 ;
      RECT  531.38 4.16 534.92 7.1 ;
      RECT  531.38 7.1 534.92 121.12 ;
      RECT  1.66 391.98 4.16 418.28 ;
      RECT  1.66 418.28 4.16 421.22 ;
      RECT  4.16 391.98 531.38 418.28 ;
      RECT  531.38 391.98 533.88 418.28 ;
      RECT  531.38 418.28 533.88 421.22 ;
      RECT  0.62 164.86 0.76 421.68 ;
      RECT  0.62 421.68 0.76 424.62 ;
      RECT  0.62 424.62 0.76 424.76 ;
      RECT  0.76 164.86 1.66 421.68 ;
      RECT  0.76 424.62 1.66 424.76 ;
      RECT  533.88 391.98 534.78 421.68 ;
      RECT  533.88 424.62 534.78 424.76 ;
      RECT  534.78 391.98 534.92 421.68 ;
      RECT  534.78 421.68 534.92 424.62 ;
      RECT  534.78 424.62 534.92 424.76 ;
      RECT  1.66 421.22 4.16 421.68 ;
      RECT  1.66 424.62 4.16 424.76 ;
      RECT  4.16 421.22 531.38 421.68 ;
      RECT  4.16 424.62 531.38 424.76 ;
      RECT  531.38 421.22 533.88 421.68 ;
      RECT  531.38 424.62 533.88 424.76 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 3.7 ;
      RECT  0.62 3.7 0.76 20.48 ;
      RECT  0.76 0.62 1.66 0.76 ;
      RECT  0.76 3.7 1.66 20.48 ;
      RECT  1.66 0.62 4.16 0.76 ;
      RECT  1.66 3.7 4.16 4.16 ;
      RECT  4.16 0.62 531.38 0.76 ;
      RECT  4.16 3.7 531.38 4.16 ;
      RECT  531.38 0.62 534.78 0.76 ;
      RECT  531.38 3.7 534.78 4.16 ;
      RECT  534.78 0.62 534.92 0.76 ;
      RECT  534.78 0.76 534.92 3.7 ;
      RECT  534.78 3.7 534.92 4.16 ;
   LAYER  met4 ;
      RECT  105.7 0.62 110.24 1.66 ;
      RECT  111.82 0.62 115.68 1.66 ;
      RECT  117.26 0.62 122.48 1.66 ;
      RECT  124.06 0.62 127.92 1.66 ;
      RECT  129.5 0.62 133.36 1.66 ;
      RECT  134.94 0.62 139.48 1.66 ;
      RECT  141.06 0.62 144.92 1.66 ;
      RECT  146.5 0.62 151.72 1.66 ;
      RECT  153.3 0.62 157.16 1.66 ;
      RECT  158.74 0.62 162.6 1.66 ;
      RECT  363.42 0.62 367.28 1.66 ;
      RECT  374.3 0.62 378.84 1.66 ;
      RECT  380.42 0.62 384.28 1.66 ;
      RECT  385.86 0.62 391.08 1.66 ;
      RECT  392.66 0.62 396.52 1.66 ;
      RECT  398.1 0.62 401.96 1.66 ;
      RECT  403.54 0.62 408.76 1.66 ;
      RECT  410.34 0.62 414.2 1.66 ;
      RECT  415.78 0.62 419.64 1.66 ;
      RECT  421.22 0.62 425.76 1.66 ;
      RECT  427.34 0.62 431.2 1.66 ;
      RECT  450.46 0.62 454.32 1.66 ;
      RECT  455.9 0.62 460.44 1.66 ;
      RECT  462.02 0.62 466.56 1.66 ;
      RECT  468.14 0.62 472.68 1.66 ;
      RECT  51.08 1.66 52.66 423.72 ;
      RECT  52.66 1.66 104.12 423.72 ;
      RECT  52.66 423.72 57.88 424.76 ;
      RECT  59.46 423.72 64.0 424.76 ;
      RECT  65.58 423.72 69.44 424.76 ;
      RECT  71.02 423.72 74.88 424.76 ;
      RECT  76.46 423.72 80.32 424.76 ;
      RECT  81.9 423.72 87.12 424.76 ;
      RECT  88.7 423.72 92.56 424.76 ;
      RECT  94.14 423.72 98.0 424.76 ;
      RECT  99.58 423.72 104.12 424.76 ;
      RECT  104.12 1.66 104.8 423.72 ;
      RECT  104.12 423.72 104.8 424.76 ;
      RECT  104.8 1.66 105.7 423.72 ;
      RECT  105.7 1.66 106.38 423.72 ;
      RECT  106.38 423.72 110.24 424.76 ;
      RECT  111.82 423.72 116.36 424.76 ;
      RECT  117.94 423.72 121.8 424.76 ;
      RECT  123.38 423.72 127.24 424.76 ;
      RECT  128.82 423.72 133.36 424.76 ;
      RECT  134.94 423.72 139.48 424.76 ;
      RECT  141.06 423.72 145.6 424.76 ;
      RECT  147.18 423.72 151.04 424.76 ;
      RECT  152.62 423.72 156.48 424.76 ;
      RECT  158.06 423.72 162.6 424.76 ;
      RECT  374.98 423.72 378.84 424.76 ;
      RECT  380.42 423.72 384.96 424.76 ;
      RECT  386.54 423.72 390.4 424.76 ;
      RECT  391.98 423.72 395.84 424.76 ;
      RECT  397.42 423.72 401.96 424.76 ;
      RECT  403.54 423.72 408.08 424.76 ;
      RECT  409.66 423.72 413.52 424.76 ;
      RECT  415.1 423.72 418.96 424.76 ;
      RECT  432.78 0.62 437.32 1.66 ;
      RECT  445.7 0.62 448.88 1.66 ;
      RECT  442.98 0.62 443.44 1.66 ;
      RECT  31.58 0.62 104.12 1.66 ;
      RECT  164.18 0.62 166.68 1.66 ;
      RECT  168.26 0.62 168.72 1.66 ;
      RECT  170.3 0.62 172.12 1.66 ;
      RECT  174.38 0.62 174.84 1.66 ;
      RECT  176.42 0.62 178.24 1.66 ;
      RECT  179.82 0.62 180.28 1.66 ;
      RECT  183.22 0.62 184.36 1.66 ;
      RECT  187.98 0.62 191.84 1.66 ;
      RECT  194.78 0.62 197.96 1.66 ;
      RECT  200.9 0.62 203.4 1.66 ;
      RECT  206.34 0.62 209.52 1.66 ;
      RECT  212.46 0.62 214.96 1.66 ;
      RECT  218.58 0.62 221.08 1.66 ;
      RECT  225.38 0.62 227.2 1.66 ;
      RECT  228.78 0.62 229.24 1.66 ;
      RECT  231.5 0.62 233.32 1.66 ;
      RECT  237.62 0.62 238.76 1.66 ;
      RECT  240.34 0.62 240.8 1.66 ;
      RECT  243.74 0.62 244.2 1.66 ;
      RECT  245.78 0.62 247.6 1.66 ;
      RECT  249.86 0.62 251.0 1.66 ;
      RECT  252.58 0.62 253.72 1.66 ;
      RECT  255.98 0.62 256.44 1.66 ;
      RECT  258.02 0.62 259.84 1.66 ;
      RECT  261.42 0.62 261.88 1.66 ;
      RECT  264.82 0.62 265.96 1.66 ;
      RECT  267.54 0.62 268.0 1.66 ;
      RECT  270.26 0.62 272.08 1.66 ;
      RECT  275.7 0.62 277.52 1.66 ;
      RECT  279.1 0.62 279.56 1.66 ;
      RECT  281.82 0.62 283.64 1.66 ;
      RECT  285.22 0.62 285.68 1.66 ;
      RECT  287.94 0.62 291.12 1.66 ;
      RECT  294.06 0.62 297.24 1.66 ;
      RECT  300.18 0.62 302.68 1.66 ;
      RECT  306.3 0.62 309.48 1.66 ;
      RECT  312.42 0.62 314.92 1.66 ;
      RECT  318.54 0.62 320.36 1.66 ;
      RECT  321.94 0.62 322.4 1.66 ;
      RECT  324.66 0.62 327.16 1.66 ;
      RECT  331.46 0.62 332.6 1.66 ;
      RECT  334.18 0.62 334.64 1.66 ;
      RECT  337.58 0.62 338.04 1.66 ;
      RECT  339.62 0.62 340.76 1.66 ;
      RECT  345.06 0.62 347.56 1.66 ;
      RECT  349.14 0.62 349.6 1.66 ;
      RECT  351.86 0.62 353.0 1.66 ;
      RECT  356.62 0.62 359.12 1.66 ;
      RECT  360.7 0.62 361.16 1.66 ;
      RECT  369.54 0.62 372.72 1.66 ;
      RECT  164.18 423.72 166.0 424.76 ;
      RECT  167.58 423.72 168.72 424.76 ;
      RECT  170.3 423.72 172.12 424.76 ;
      RECT  173.7 423.72 174.16 424.76 ;
      RECT  177.1 423.72 178.24 424.76 ;
      RECT  181.18 423.72 181.64 424.76 ;
      RECT  183.22 423.72 185.72 424.76 ;
      RECT  188.66 423.72 191.84 424.76 ;
      RECT  194.78 423.72 197.28 424.76 ;
      RECT  200.22 423.72 203.4 424.76 ;
      RECT  206.34 423.72 208.84 424.76 ;
      RECT  212.46 423.72 215.64 424.76 ;
      RECT  218.58 423.72 221.08 424.76 ;
      RECT  225.38 423.72 227.2 424.76 ;
      RECT  228.78 423.72 229.24 424.76 ;
      RECT  231.5 423.72 231.96 424.76 ;
      RECT  233.54 423.72 234.68 424.76 ;
      RECT  237.62 423.72 238.08 424.76 ;
      RECT  239.66 423.72 240.8 424.76 ;
      RECT  243.74 423.72 244.88 424.76 ;
      RECT  246.46 423.72 247.6 424.76 ;
      RECT  249.86 423.72 250.32 424.76 ;
      RECT  251.9 423.72 253.72 424.76 ;
      RECT  255.3 423.72 255.76 424.76 ;
      RECT  258.02 423.72 259.84 424.76 ;
      RECT  262.78 423.72 263.24 424.76 ;
      RECT  264.82 423.72 267.32 424.76 ;
      RECT  270.94 423.72 273.44 424.76 ;
      RECT  277.06 423.72 277.52 424.76 ;
      RECT  279.1 423.72 279.56 424.76 ;
      RECT  281.82 423.72 285.0 424.76 ;
      RECT  287.94 423.72 290.44 424.76 ;
      RECT  294.06 423.72 297.24 424.76 ;
      RECT  300.18 423.72 303.36 424.76 ;
      RECT  306.3 423.72 308.8 424.76 ;
      RECT  312.42 423.72 314.24 424.76 ;
      RECT  315.82 423.72 316.28 424.76 ;
      RECT  318.54 423.72 319.68 424.76 ;
      RECT  321.26 423.72 322.4 424.76 ;
      RECT  324.66 423.72 326.48 424.76 ;
      RECT  328.06 423.72 328.52 424.76 ;
      RECT  331.46 423.72 331.92 424.76 ;
      RECT  333.5 423.72 334.64 424.76 ;
      RECT  336.9 423.72 337.36 424.76 ;
      RECT  338.94 423.72 340.76 424.76 ;
      RECT  343.02 423.72 344.16 424.76 ;
      RECT  345.74 423.72 347.56 424.76 ;
      RECT  349.14 423.72 349.6 424.76 ;
      RECT  351.86 423.72 353.0 424.76 ;
      RECT  354.58 423.72 355.72 424.76 ;
      RECT  357.98 423.72 359.12 424.76 ;
      RECT  362.74 423.72 366.6 424.76 ;
      RECT  368.86 423.72 373.4 424.76 ;
      RECT  4.16 1.66 7.1 4.16 ;
      RECT  4.16 421.22 7.1 423.72 ;
      RECT  7.1 1.66 51.08 4.16 ;
      RECT  7.1 4.16 51.08 421.22 ;
      RECT  7.1 421.22 51.08 423.72 ;
      RECT  106.38 1.66 528.44 4.16 ;
      RECT  106.38 4.16 528.44 421.22 ;
      RECT  106.38 421.22 528.44 423.72 ;
      RECT  528.44 1.66 531.38 4.16 ;
      RECT  528.44 421.22 531.38 423.72 ;
      RECT  474.26 0.62 531.84 0.76 ;
      RECT  474.26 0.76 531.84 1.66 ;
      RECT  531.84 0.62 534.78 0.76 ;
      RECT  534.78 0.62 534.92 0.76 ;
      RECT  534.78 0.76 534.92 1.66 ;
      RECT  420.54 423.72 531.84 424.62 ;
      RECT  420.54 424.62 531.84 424.76 ;
      RECT  531.84 424.62 534.78 424.76 ;
      RECT  534.78 423.72 534.92 424.62 ;
      RECT  534.78 424.62 534.92 424.76 ;
      RECT  531.38 1.66 531.84 4.16 ;
      RECT  534.78 1.66 534.92 4.16 ;
      RECT  531.38 4.16 531.84 421.22 ;
      RECT  534.78 4.16 534.92 421.22 ;
      RECT  531.38 421.22 531.84 423.72 ;
      RECT  534.78 421.22 534.92 423.72 ;
      RECT  0.62 423.72 0.76 424.62 ;
      RECT  0.62 424.62 0.76 424.76 ;
      RECT  0.76 424.62 3.7 424.76 ;
      RECT  3.7 423.72 51.08 424.62 ;
      RECT  3.7 424.62 51.08 424.76 ;
      RECT  0.62 0.62 0.76 0.76 ;
      RECT  0.62 0.76 0.76 1.66 ;
      RECT  0.76 0.62 3.7 0.76 ;
      RECT  3.7 0.62 30.0 0.76 ;
      RECT  3.7 0.76 30.0 1.66 ;
      RECT  0.62 1.66 0.76 4.16 ;
      RECT  3.7 1.66 4.16 4.16 ;
      RECT  0.62 4.16 0.76 421.22 ;
      RECT  3.7 4.16 4.16 421.22 ;
      RECT  0.62 421.22 0.76 423.72 ;
      RECT  3.7 421.22 4.16 423.72 ;
   END
END    sky130_sram_2rw_64x128_64
END    LIBRARY
